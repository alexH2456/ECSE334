* C:\Users\zizou\ECSE334\Assignment3\Draft2.asc
M1 N002 N005 N007 N007 QMOS1
M2 N001 N006 N007 N007 QMOS1
M5 N001 N003 N006 N006 QMOS1

I1 N007 N004 200uA
I3 N006 N004 0.8mA
I2 N003 N004 300uA

M4 N003 N002 N001 N001 QMOS4
M3 N002 N002 N001 N001 QMOS3

VS N005 0 AC 1
VSS N004 0 -2.5V
VDD N001 0 +2.5V

.model QMOS1 NMOS (LEVEL=2 L=1u W=20u VTo=0.7 Kp=0.12m LAMBDA=41.66667m)
.model QMOS3 PMOS (LEVEL=2 L=1u W=40u VTo=-0.7 Kp=0.06m LAMBDA=41.66667m)
.model QMOS4 PMOS (LEVEL=2 L=1u W=120u VTo=-0.7 Kp=0.06m LAMBDA=41.66667m)
.lib E:\My Documents\LTspiceXVII\lib\cmp\standard.mos
.backanno

.op
.ac dec 100 1 10k

.end
