ECSE 334 - Assignment 3

*Voltage Sources
Vs g1 0 0V
Vcc s3 0 2.5V
Vss i1 0 -2.5V

*Current Sources
I1 s1 i1 200uA
I2 op i1 0.8mA
I3 g5 i1 300uA

*PMOS Transistors
M4 g5 d1 s3 p QMOS4
M3 d1 d1 s3 p QMOS3

*NMOS Transistors
M1 d1 g1 s1 n QMOS125
M2 s3 op s1 n QMOS125
M5 s3 g5 op n QMOS125

.model QMOS3 PMOS(LEVEL=2 L=1 W=40 VTo=-0.7 Kp=0.06m LAMBDA=0.0417)
.model QMOS4 PMOS(LEVEL=2 L=1 W=120 VTo=-0.7 Kp=0.06m LAMBDA=0.0417)
.model QMOS125 NMOS(LEVEL=2 L=1 W=20 VTo=0.7 Kp=0.12m LAMBDA=0.0417)

.op

.end
