Assignment 1

*Voltage Sources
VCC 3 0 5V

*PNP Transistors
Q1 b b 3 QPNP
Q2 rl b 3 QPNP

*Design Param
Ref b 0 1kohm
Rl rl 0 1kohm


.model QPNP	PNP (Is=1f Xti=3 Eg=1.11 Vaf=50 Bf=50 Ne=1.5 Ise=0 Ikf=80m Xtb=1.5 Br=4.977 Nc=2 Isc=0 Ikr=0 Rc=2.5 Cjc=9.728p Mjc=.5776 Vjc=.75 Fc=.5 Cje=8.063p Mje=.3677 Vje=.75 Tr=33.42n Tf=179.3p Itf=.4 Vtf=4 Xtf=6 Rb=10)
*		National	pid=66		case=TO92
*		88-09-09 bam	creation

.OP

.END
